mem['h0000] = 32'h00000517;
mem['h0001] = 32'h66850513;
mem['h0002] = 32'h10000597;
mem['h0003] = 32'hFF858593;
mem['h0004] = 32'h10000617;
mem['h0005] = 32'hFF060613;
mem['h0006] = 32'h00C5DC63;
mem['h0007] = 32'h00052683;
mem['h0008] = 32'h00D5A023;
mem['h0009] = 32'h00450513;
mem['h000A] = 32'h00458593;
mem['h000B] = 32'hFEC5C8E3;
mem['h000C] = 32'h10000517;
mem['h000D] = 32'hFD050513;
mem['h000E] = 32'h00418593;
mem['h000F] = 32'h00B55863;
mem['h0010] = 32'h00052023;
mem['h0011] = 32'h00450513;
mem['h0012] = 32'hFEB54CE3;
mem['h0013] = 32'h10008117;
mem['h0014] = 32'hFB410113;
mem['h0015] = 32'h10000197;
mem['h0016] = 32'h7AC18193;
mem['h0017] = 32'h00A54533;
mem['h0018] = 32'h00B5C5B3;
mem['h0019] = 32'h00C64633;
mem['h001A] = 32'h1BC000EF;
mem['h001B] = 32'h0000006F;
mem['h001C] = 32'h00052783;
mem['h001D] = 32'h0087A783;
mem['h001E] = 32'h0007A783;
mem['h001F] = 32'h0007A783;
mem['h0020] = 32'hFE07C8E3;
mem['h0021] = 32'h00052783;
mem['h0022] = 32'h0087A783;
mem['h0023] = 32'h0007A783;
mem['h0024] = 32'h00B78023;
mem['h0025] = 32'h00008067;
mem['h0026] = 32'h0A058A63;
mem['h0027] = 32'hFE010113;
mem['h0028] = 32'h00912A23;
mem['h0029] = 32'h00058493;
mem['h002A] = 32'h01212823;
mem['h002B] = 32'h00A00593;
mem['h002C] = 32'h00050913;
mem['h002D] = 32'h00048513;
mem['h002E] = 32'h00812C23;
mem['h002F] = 32'h00112E23;
mem['h0030] = 32'h01312623;
mem['h0031] = 32'h01412423;
mem['h0032] = 32'h4A4000EF;
mem['h0033] = 32'h01051513;
mem['h0034] = 32'h01055513;
mem['h0035] = 32'h00100413;
mem['h0036] = 32'h06857E63;
mem['h0037] = 32'h00900A13;
mem['h0038] = 32'h00040593;
mem['h0039] = 32'h00048513;
mem['h003A] = 32'h484000EF;
mem['h003B] = 32'h03050593;
mem['h003C] = 32'h0FF5F593;
mem['h003D] = 32'h00090513;
mem['h003E] = 32'hF79FF0EF;
mem['h003F] = 32'h00040593;
mem['h0040] = 32'h00048513;
mem['h0041] = 32'h4B0000EF;
mem['h0042] = 32'h01051493;
mem['h0043] = 32'h00A00593;
mem['h0044] = 32'h00040513;
mem['h0045] = 32'h458000EF;
mem['h0046] = 32'h00040993;
mem['h0047] = 32'h01051413;
mem['h0048] = 32'h0104D493;
mem['h0049] = 32'h01045413;
mem['h004A] = 32'hFB3A6CE3;
mem['h004B] = 32'h01C12083;
mem['h004C] = 32'h01812403;
mem['h004D] = 32'h01412483;
mem['h004E] = 32'h01012903;
mem['h004F] = 32'h00C12983;
mem['h0050] = 32'h00812A03;
mem['h0051] = 32'h02010113;
mem['h0052] = 32'h00008067;
mem['h0053] = 32'h03000593;
mem['h0054] = 32'hF21FF06F;
mem['h0055] = 32'h00241793;
mem['h0056] = 32'h00F40433;
mem['h0057] = 32'h00141413;
mem['h0058] = 32'h01041413;
mem['h0059] = 32'h01045413;
mem['h005A] = 32'hF71FF06F;
mem['h005B] = 32'hFF010113;
mem['h005C] = 32'h00812423;
mem['h005D] = 32'h00912223;
mem['h005E] = 32'h00112623;
mem['h005F] = 32'h00050493;
mem['h0060] = 32'h00058413;
mem['h0061] = 32'h00044583;
mem['h0062] = 32'h00059C63;
mem['h0063] = 32'h00C12083;
mem['h0064] = 32'h00812403;
mem['h0065] = 32'h00412483;
mem['h0066] = 32'h01010113;
mem['h0067] = 32'h00008067;
mem['h0068] = 32'h00048513;
mem['h0069] = 32'h00140413;
mem['h006A] = 32'hEC9FF0EF;
mem['h006B] = 32'hFD9FF06F;
mem['h006C] = 32'h0001A703;
mem['h006D] = 32'h100007B7;
mem['h006E] = 32'h00078793;
mem['h006F] = 32'h00F707B3;
mem['h0070] = 32'h00A70733;
mem['h0071] = 32'h00E1A023;
mem['h0072] = 32'h000016B7;
mem['h0073] = 32'h80068693;
mem['h0074] = 32'h00E6D463;
mem['h0075] = 32'h00100073;
mem['h0076] = 32'h00078513;
mem['h0077] = 32'h00008067;
mem['h0078] = 32'h0FF5F593;
mem['h0079] = 32'h00000793;
mem['h007A] = 32'h00C79463;
mem['h007B] = 32'h00008067;
mem['h007C] = 32'h00F50733;
mem['h007D] = 32'h00B70023;
mem['h007E] = 32'h00178793;
mem['h007F] = 32'hFEDFF06F;
mem['h0080] = 32'h00000793;
mem['h0081] = 32'h00C79463;
mem['h0082] = 32'h00008067;
mem['h0083] = 32'h00F58733;
mem['h0084] = 32'h00074683;
mem['h0085] = 32'h00F50733;
mem['h0086] = 32'h00178793;
mem['h0087] = 32'h00D70023;
mem['h0088] = 32'hFE5FF06F;
mem['h0089] = 32'hFB010113;
mem['h008A] = 32'h01000513;
mem['h008B] = 32'h04112623;
mem['h008C] = 32'h04812423;
mem['h008D] = 32'h04912223;
mem['h008E] = 32'h03312E23;
mem['h008F] = 32'h03412C23;
mem['h0090] = 32'h03512A23;
mem['h0091] = 32'h03612823;
mem['h0092] = 32'h05212023;
mem['h0093] = 32'h03712623;
mem['h0094] = 32'h03812423;
mem['h0095] = 32'hF5DFF0EF;
mem['h0096] = 32'h00050413;
mem['h0097] = 32'h01000513;
mem['h0098] = 32'hF51FF0EF;
mem['h0099] = 32'h00050493;
mem['h009A] = 32'h00400513;
mem['h009B] = 32'hF45FF0EF;
mem['h009C] = 32'h200007B7;
mem['h009D] = 32'h00F52023;
mem['h009E] = 32'h00A4A023;
mem['h009F] = 32'h00400513;
mem['h00A0] = 32'hF31FF0EF;
mem['h00A1] = 32'h200007B7;
mem['h00A2] = 32'h00478793;
mem['h00A3] = 32'h00F52023;
mem['h00A4] = 32'h00A4A223;
mem['h00A5] = 32'h00400513;
mem['h00A6] = 32'hF19FF0EF;
mem['h00A7] = 32'h200007B7;
mem['h00A8] = 32'h00878793;
mem['h00A9] = 32'h00F52023;
mem['h00AA] = 32'h00A4A423;
mem['h00AB] = 32'h00400513;
mem['h00AC] = 32'hF01FF0EF;
mem['h00AD] = 32'h200007B7;
mem['h00AE] = 32'h00C78793;
mem['h00AF] = 32'h00F52023;
mem['h00B0] = 32'h00A4A623;
mem['h00B1] = 32'h00942023;
mem['h00B2] = 32'h00400513;
mem['h00B3] = 32'hEE5FF0EF;
mem['h00B4] = 32'h200007B7;
mem['h00B5] = 32'h01078793;
mem['h00B6] = 32'h00F52023;
mem['h00B7] = 32'h00A42223;
mem['h00B8] = 32'h00400513;
mem['h00B9] = 32'hECDFF0EF;
mem['h00BA] = 32'h200007B7;
mem['h00BB] = 32'h01478793;
mem['h00BC] = 32'h00F52023;
mem['h00BD] = 32'h00A42423;
mem['h00BE] = 32'h00400513;
mem['h00BF] = 32'hEB5FF0EF;
mem['h00C0] = 32'h200007B7;
mem['h00C1] = 32'h01878793;
mem['h00C2] = 32'h00F52023;
mem['h00C3] = 32'h00442783;
mem['h00C4] = 32'h00A42623;
mem['h00C5] = 32'h0007A703;
mem['h00C6] = 32'h61800593;
mem['h00C7] = 32'h00040513;
mem['h00C8] = 32'h00072783;
mem['h00C9] = 32'h01200A93;
mem['h00CA] = 32'h00A00993;
mem['h00CB] = 32'h2007E793;
mem['h00CC] = 32'h00F72023;
mem['h00CD] = 32'h00442703;
mem['h00CE] = 32'h00442783;
mem['h00CF] = 32'h00D00A13;
mem['h00D0] = 32'h00072683;
mem['h00D1] = 32'h0007A783;
mem['h00D2] = 32'h07F00B13;
mem['h00D3] = 32'h0007A703;
mem['h00D4] = 32'h0006A783;
mem['h00D5] = 32'h00177713;
mem['h00D6] = 32'h00871713;
mem['h00D7] = 32'hEFF7F793;
mem['h00D8] = 32'h00E7E7B3;
mem['h00D9] = 32'h00F6A023;
mem['h00DA] = 32'hE05FF0EF;
mem['h00DB] = 32'h00042783;
mem['h00DC] = 32'h0007A783;
mem['h00DD] = 32'h0007A783;
mem['h00DE] = 32'h0007A583;
mem['h00DF] = 32'hFE05D8E3;
mem['h00E0] = 32'h0FF5F793;
mem['h00E1] = 32'hFF5784E3;
mem['h00E2] = 32'h0FF5F593;
mem['h00E3] = 32'h00B10023;
mem['h00E4] = 32'hFD358EE3;
mem['h00E5] = 32'h00000493;
mem['h00E6] = 32'h00010913;
mem['h00E7] = 32'h07458663;
mem['h00E8] = 32'h00800C13;
mem['h00E9] = 32'h01F00B93;
mem['h00EA] = 32'h01858463;
mem['h00EB] = 32'h1B659263;
mem['h00EC] = 32'h02905863;
mem['h00ED] = 32'h00800593;
mem['h00EE] = 32'h00040513;
mem['h00EF] = 32'hCB5FF0EF;
mem['h00F0] = 32'h02000593;
mem['h00F1] = 32'h00040513;
mem['h00F2] = 32'hCA9FF0EF;
mem['h00F3] = 32'h00800593;
mem['h00F4] = 32'h00040513;
mem['h00F5] = 32'hFFF90913;
mem['h00F6] = 32'hFFF48493;
mem['h00F7] = 32'hC95FF0EF;
mem['h00F8] = 32'h00042783;
mem['h00F9] = 32'h0007A783;
mem['h00FA] = 32'h0007A783;
mem['h00FB] = 32'h0007A583;
mem['h00FC] = 32'hFE05D8E3;
mem['h00FD] = 32'h03748663;
mem['h00FE] = 32'h0FF5F593;
mem['h00FF] = 32'h00B90023;
mem['h0100] = 32'h03358063;
mem['h0101] = 32'hFB4592E3;
mem['h0102] = 32'h00D00593;
mem['h0103] = 32'h00040513;
mem['h0104] = 32'hC61FF0EF;
mem['h0105] = 32'h00A00593;
mem['h0106] = 32'h00040513;
mem['h0107] = 32'hC55FF0EF;
mem['h0108] = 32'h00090023;
mem['h0109] = 32'h0FF4F493;
mem['h010A] = 32'hF40482E3;
mem['h010B] = 32'h62800593;
mem['h010C] = 32'h00040513;
mem['h010D] = 32'hD39FF0EF;
mem['h010E] = 32'h00842783;
mem['h010F] = 32'h00C00493;
mem['h0110] = 32'h0007A783;
mem['h0111] = 32'h65400913;
mem['h0112] = 32'hFFC00993;
mem['h0113] = 32'h0027DA03;
mem['h0114] = 32'h009A57B3;
mem['h0115] = 32'h00F7F793;
mem['h0116] = 32'h00F907B3;
mem['h0117] = 32'h0007C583;
mem['h0118] = 32'h00040513;
mem['h0119] = 32'hFFC48493;
mem['h011A] = 32'hC09FF0EF;
mem['h011B] = 32'hFF3492E3;
mem['h011C] = 32'h63400593;
mem['h011D] = 32'h00040513;
mem['h011E] = 32'hCF5FF0EF;
mem['h011F] = 32'h00842783;
mem['h0120] = 32'h00C00493;
mem['h0121] = 32'hFFC00993;
mem['h0122] = 32'h0007A783;
mem['h0123] = 32'h0007DA03;
mem['h0124] = 32'h009A57B3;
mem['h0125] = 32'h00F7F793;
mem['h0126] = 32'h00F907B3;
mem['h0127] = 32'h0007C583;
mem['h0128] = 32'h00040513;
mem['h0129] = 32'hFFC48493;
mem['h012A] = 32'hBC9FF0EF;
mem['h012B] = 32'hFF3492E3;
mem['h012C] = 32'h00040513;
mem['h012D] = 32'h64400593;
mem['h012E] = 32'hCB5FF0EF;
mem['h012F] = 32'h00C42783;
mem['h0130] = 32'h00040513;
mem['h0131] = 32'h0007A783;
mem['h0132] = 32'h0037C583;
mem['h0133] = 32'hBCDFF0EF;
mem['h0134] = 32'h00040513;
mem['h0135] = 32'h02E00593;
mem['h0136] = 32'hB99FF0EF;
mem['h0137] = 32'h00C42783;
mem['h0138] = 32'h00040513;
mem['h0139] = 32'h0007A783;
mem['h013A] = 32'h0027C583;
mem['h013B] = 32'hBADFF0EF;
mem['h013C] = 32'h00040513;
mem['h013D] = 32'h02E00593;
mem['h013E] = 32'hB79FF0EF;
mem['h013F] = 32'h00C42783;
mem['h0140] = 32'h00040513;
mem['h0141] = 32'h0007A783;
mem['h0142] = 32'h0007D583;
mem['h0143] = 32'hB8DFF0EF;
mem['h0144] = 32'h00040513;
mem['h0145] = 32'h62400593;
mem['h0146] = 32'hC55FF0EF;
mem['h0147] = 32'h04C12083;
mem['h0148] = 32'h04812403;
mem['h0149] = 32'h04412483;
mem['h014A] = 32'h04012903;
mem['h014B] = 32'h03C12983;
mem['h014C] = 32'h03812A03;
mem['h014D] = 32'h03412A83;
mem['h014E] = 32'h03012B03;
mem['h014F] = 32'h02C12B83;
mem['h0150] = 32'h02812C03;
mem['h0151] = 32'h00000513;
mem['h0152] = 32'h05010113;
mem['h0153] = 32'h00008067;
mem['h0154] = 32'h00040513;
mem['h0155] = 32'hB1DFF0EF;
mem['h0156] = 32'h00190913;
mem['h0157] = 32'h00148493;
mem['h0158] = 32'hE81FF06F;
mem['h0159] = 32'h06054063;
mem['h015A] = 32'h0605C663;
mem['h015B] = 32'h00058613;
mem['h015C] = 32'h00050593;
mem['h015D] = 32'hFFF00513;
mem['h015E] = 32'h02060C63;
mem['h015F] = 32'h00100693;
mem['h0160] = 32'h00B67A63;
mem['h0161] = 32'h00C05863;
mem['h0162] = 32'h00161613;
mem['h0163] = 32'h00169693;
mem['h0164] = 32'hFEB66AE3;
mem['h0165] = 32'h00000513;
mem['h0166] = 32'h00C5E663;
mem['h0167] = 32'h40C585B3;
mem['h0168] = 32'h00D56533;
mem['h0169] = 32'h0016D693;
mem['h016A] = 32'h00165613;
mem['h016B] = 32'hFE0696E3;
mem['h016C] = 32'h00008067;
mem['h016D] = 32'h00008293;
mem['h016E] = 32'hFB5FF0EF;
mem['h016F] = 32'h00058513;
mem['h0170] = 32'h00028067;
mem['h0171] = 32'h40A00533;
mem['h0172] = 32'h00B04863;
mem['h0173] = 32'h40B005B3;
mem['h0174] = 32'hF9DFF06F;
mem['h0175] = 32'h40B005B3;
mem['h0176] = 32'h00008293;
mem['h0177] = 32'hF91FF0EF;
mem['h0178] = 32'h40A00533;
mem['h0179] = 32'h00028067;
mem['h017A] = 32'h00008293;
mem['h017B] = 32'h0005CA63;
mem['h017C] = 32'h00054C63;
mem['h017D] = 32'hF79FF0EF;
mem['h017E] = 32'h00058513;
mem['h017F] = 32'h00028067;
mem['h0180] = 32'h40B005B3;
mem['h0181] = 32'hFE0558E3;
mem['h0182] = 32'h40A00533;
mem['h0183] = 32'hF61FF0EF;
mem['h0184] = 32'h40B00533;
mem['h0185] = 32'h00028067;
mem['h0186] = 32'h6C6C6548;
mem['h0187] = 32'h6F77206F;
mem['h0188] = 32'h21646C72;
mem['h0189] = 32'h00000A0D;
mem['h018A] = 32'h444E4556;
mem['h018B] = 32'h2020524F;
mem['h018C] = 32'h0000203D;
mem['h018D] = 32'h52500A0D;
mem['h018E] = 32'h4355444F;
mem['h018F] = 32'h203D2054;
mem['h0190] = 32'h00000000;
mem['h0191] = 32'h45560A0D;
mem['h0192] = 32'h4F495352;
mem['h0193] = 32'h203D204E;
mem['h0194] = 32'h00000076;
mem['h0195] = 32'h33323130;
mem['h0196] = 32'h37363534;
mem['h0197] = 32'h42413938;
mem['h0198] = 32'h46454443;
mem['h0199] = 32'h00000000;
