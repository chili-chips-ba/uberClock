mem['h0000] = 32'h00000517;
mem['h0001] = 32'h26C50513;
mem['h0002] = 32'h10000597;
mem['h0003] = 32'hFF858593;
mem['h0004] = 32'h10000617;
mem['h0005] = 32'hFF060613;
mem['h0006] = 32'h00C5DC63;
mem['h0007] = 32'h00052683;
mem['h0008] = 32'h00D5A023;
mem['h0009] = 32'h00450513;
mem['h000A] = 32'h00458593;
mem['h000B] = 32'hFEC5C8E3;
mem['h000C] = 32'h10000517;
mem['h000D] = 32'hFD050513;
mem['h000E] = 32'h00418593;
mem['h000F] = 32'h00B55863;
mem['h0010] = 32'h00052023;
mem['h0011] = 32'h00450513;
mem['h0012] = 32'hFEB54CE3;
mem['h0013] = 32'h10008117;
mem['h0014] = 32'hFB410113;
mem['h0015] = 32'h10000197;
mem['h0016] = 32'h7AC18193;
mem['h0017] = 32'h00A54533;
mem['h0018] = 32'h00B5C5B3;
mem['h0019] = 32'h00C64633;
mem['h001A] = 32'h07C000EF;
mem['h001B] = 32'h0000006F;
mem['h001C] = 32'h0001A703;
mem['h001D] = 32'h100007B7;
mem['h001E] = 32'h00078793;
mem['h001F] = 32'h00F707B3;
mem['h0020] = 32'h00A70733;
mem['h0021] = 32'h00E1A023;
mem['h0022] = 32'h000016B7;
mem['h0023] = 32'h80068693;
mem['h0024] = 32'h00E6D463;
mem['h0025] = 32'h00100073;
mem['h0026] = 32'h00078513;
mem['h0027] = 32'h00008067;
mem['h0028] = 32'h0FF5F593;
mem['h0029] = 32'h00000793;
mem['h002A] = 32'h00C79463;
mem['h002B] = 32'h00008067;
mem['h002C] = 32'h00F50733;
mem['h002D] = 32'h00B70023;
mem['h002E] = 32'h00178793;
mem['h002F] = 32'hFEDFF06F;
mem['h0030] = 32'h00000793;
mem['h0031] = 32'h00C79463;
mem['h0032] = 32'h00008067;
mem['h0033] = 32'h00F58733;
mem['h0034] = 32'h00074683;
mem['h0035] = 32'h00F50733;
mem['h0036] = 32'h00178793;
mem['h0037] = 32'h00D70023;
mem['h0038] = 32'hFE5FF06F;
mem['h0039] = 32'hFF010113;
mem['h003A] = 32'h01800513;
mem['h003B] = 32'h00112623;
mem['h003C] = 32'h00812423;
mem['h003D] = 32'h00912223;
mem['h003E] = 32'hF79FF0EF;
mem['h003F] = 32'h00050413;
mem['h0040] = 32'h01000513;
mem['h0041] = 32'hF6DFF0EF;
mem['h0042] = 32'h00050493;
mem['h0043] = 32'h00400513;
mem['h0044] = 32'hF61FF0EF;
mem['h0045] = 32'h200007B7;
mem['h0046] = 32'h00F52023;
mem['h0047] = 32'h00A4A023;
mem['h0048] = 32'h00400513;
mem['h0049] = 32'hF4DFF0EF;
mem['h004A] = 32'h200007B7;
mem['h004B] = 32'h00478793;
mem['h004C] = 32'h00F52023;
mem['h004D] = 32'h00A4A223;
mem['h004E] = 32'h00400513;
mem['h004F] = 32'hF35FF0EF;
mem['h0050] = 32'h200007B7;
mem['h0051] = 32'h00878793;
mem['h0052] = 32'h00F52023;
mem['h0053] = 32'h00A4A423;
mem['h0054] = 32'h00400513;
mem['h0055] = 32'hF1DFF0EF;
mem['h0056] = 32'h200007B7;
mem['h0057] = 32'h00C78793;
mem['h0058] = 32'h00F52023;
mem['h0059] = 32'h00A4A623;
mem['h005A] = 32'h00942023;
mem['h005B] = 32'h00400513;
mem['h005C] = 32'hF01FF0EF;
mem['h005D] = 32'h200007B7;
mem['h005E] = 32'h01078793;
mem['h005F] = 32'h00F52023;
mem['h0060] = 32'h00A42223;
mem['h0061] = 32'h00400513;
mem['h0062] = 32'hEE9FF0EF;
mem['h0063] = 32'h200007B7;
mem['h0064] = 32'h01478793;
mem['h0065] = 32'h00F52023;
mem['h0066] = 32'h00A42423;
mem['h0067] = 32'h00400513;
mem['h0068] = 32'hED1FF0EF;
mem['h0069] = 32'h200007B7;
mem['h006A] = 32'h01878793;
mem['h006B] = 32'h00F52023;
mem['h006C] = 32'h00A42623;
mem['h006D] = 32'h00400513;
mem['h006E] = 32'hEB9FF0EF;
mem['h006F] = 32'h200007B7;
mem['h0070] = 32'h01C78793;
mem['h0071] = 32'h00F52023;
mem['h0072] = 32'h00A42823;
mem['h0073] = 32'h00400513;
mem['h0074] = 32'hEA1FF0EF;
mem['h0075] = 32'h25C00793;
mem['h0076] = 32'h0007C703;
mem['h0077] = 32'h04071A63;
mem['h0078] = 32'h00001637;
mem['h0079] = 32'h000046B7;
mem['h007A] = 32'hFFF60613;
mem['h007B] = 32'hFFF68693;
mem['h007C] = 32'hFFFFC537;
mem['h007D] = 32'h01042703;
mem['h007E] = 32'h00C42783;
mem['h007F] = 32'h00072583;
mem['h0080] = 32'h0007A783;
mem['h0081] = 32'h0005A703;
mem['h0082] = 32'h0007A783;
mem['h0083] = 32'h00A77733;
mem['h0084] = 32'h00C7F7B3;
mem['h0085] = 32'h01079793;
mem['h0086] = 32'h0107D793;
mem['h0087] = 32'h00279793;
mem['h0088] = 32'h00D7F7B3;
mem['h0089] = 32'h00F767B3;
mem['h008A] = 32'h00F5A023;
mem['h008B] = 32'hFC9FF06F;
mem['h008C] = 32'h00178793;
mem['h008D] = 32'h00042683;
mem['h008E] = 32'h0086A683;
mem['h008F] = 32'h0006A683;
mem['h0090] = 32'h0006A683;
mem['h0091] = 32'hFE06C8E3;
mem['h0092] = 32'h00042683;
mem['h0093] = 32'h0086A683;
mem['h0094] = 32'h0006A683;
mem['h0095] = 32'h00E68023;
mem['h0096] = 32'hF81FF06F;
mem['h0097] = 32'h6C6C6548;
mem['h0098] = 32'h6F77206F;
mem['h0099] = 32'h21646C72;
mem['h009A] = 32'h00000A0D;
