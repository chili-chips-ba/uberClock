mem['h0000] = 32'h00000517;
mem['h0001] = 32'h71850513;
mem['h0002] = 32'h10000597;
mem['h0003] = 32'hFF858593;
mem['h0004] = 32'h10000617;
mem['h0005] = 32'hFF060613;
mem['h0006] = 32'h00C5DC63;
mem['h0007] = 32'h00052683;
mem['h0008] = 32'h00D5A023;
mem['h0009] = 32'h00450513;
mem['h000A] = 32'h00458593;
mem['h000B] = 32'hFEC5C8E3;
mem['h000C] = 32'h10000517;
mem['h000D] = 32'hFD050513;
mem['h000E] = 32'h10000597;
mem['h000F] = 32'h7CC58593;
mem['h0010] = 32'h00B55863;
mem['h0011] = 32'h00052023;
mem['h0012] = 32'h00450513;
mem['h0013] = 32'hFEB54CE3;
mem['h0014] = 32'h10008117;
mem['h0015] = 32'hFB010113;
mem['h0016] = 32'h10000197;
mem['h0017] = 32'h7A818193;
mem['h0018] = 32'h00A54533;
mem['h0019] = 32'h00B5C5B3;
mem['h001A] = 32'h00C64633;
mem['h001B] = 32'h0DC000EF;
mem['h001C] = 32'h0000006F;
mem['h001D] = 32'h00052783;
mem['h001E] = 32'h0087A783;
mem['h001F] = 32'h0007A783;
mem['h0020] = 32'h0007A783;
mem['h0021] = 32'hFE07C8E3;
mem['h0022] = 32'h00052783;
mem['h0023] = 32'h0087A783;
mem['h0024] = 32'h0007A783;
mem['h0025] = 32'h00B78023;
mem['h0026] = 32'h00008067;
mem['h0027] = 32'hFE010113;
mem['h0028] = 32'h00812C23;
mem['h0029] = 32'h00112E23;
mem['h002A] = 32'h00058413;
mem['h002B] = 32'h00044583;
mem['h002C] = 32'h00059A63;
mem['h002D] = 32'h01C12083;
mem['h002E] = 32'h01812403;
mem['h002F] = 32'h02010113;
mem['h0030] = 32'h00008067;
mem['h0031] = 32'h00A12623;
mem['h0032] = 32'hFADFF0EF;
mem['h0033] = 32'h00C12503;
mem['h0034] = 32'h00140413;
mem['h0035] = 32'hFD9FF06F;
mem['h0036] = 32'h0001A703;
mem['h0037] = 32'h100007B7;
mem['h0038] = 32'h00078793;
mem['h0039] = 32'h00F707B3;
mem['h003A] = 32'h00A70733;
mem['h003B] = 32'h00E1A023;
mem['h003C] = 32'h000016B7;
mem['h003D] = 32'h80068693;
mem['h003E] = 32'h00E6D463;
mem['h003F] = 32'h00100073;
mem['h0040] = 32'h00078513;
mem['h0041] = 32'h00008067;
mem['h0042] = 32'h00000793;
mem['h0043] = 32'h00C79463;
mem['h0044] = 32'h00008067;
mem['h0045] = 32'h00F50733;
mem['h0046] = 32'h00B70023;
mem['h0047] = 32'h00178793;
mem['h0048] = 32'hFEDFF06F;
mem['h0049] = 32'h00000793;
mem['h004A] = 32'h00C79463;
mem['h004B] = 32'h00008067;
mem['h004C] = 32'h00F58733;
mem['h004D] = 32'h00074683;
mem['h004E] = 32'h00F50733;
mem['h004F] = 32'h00178793;
mem['h0050] = 32'h00D70023;
mem['h0051] = 32'hFE5FF06F;
mem['h0052] = 32'hFB010113;
mem['h0053] = 32'h01800513;
mem['h0054] = 32'h04112623;
mem['h0055] = 32'h04812423;
mem['h0056] = 32'h04912223;
mem['h0057] = 32'h05212023;
mem['h0058] = 32'h03312E23;
mem['h0059] = 32'h03412C23;
mem['h005A] = 32'h03512A23;
mem['h005B] = 32'h03612823;
mem['h005C] = 32'h03712623;
mem['h005D] = 32'h03812423;
mem['h005E] = 32'h03912223;
mem['h005F] = 32'h03A12023;
mem['h0060] = 32'h01B12E23;
mem['h0061] = 32'hF55FF0EF;
mem['h0062] = 32'h00050413;
mem['h0063] = 32'h01000513;
mem['h0064] = 32'hF49FF0EF;
mem['h0065] = 32'h00050493;
mem['h0066] = 32'h00400513;
mem['h0067] = 32'hF3DFF0EF;
mem['h0068] = 32'h200007B7;
mem['h0069] = 32'h00F52023;
mem['h006A] = 32'h00A4A023;
mem['h006B] = 32'h00400513;
mem['h006C] = 32'hF29FF0EF;
mem['h006D] = 32'h200007B7;
mem['h006E] = 32'h00478793;
mem['h006F] = 32'h00F52023;
mem['h0070] = 32'h00A4A223;
mem['h0071] = 32'h00400513;
mem['h0072] = 32'hF11FF0EF;
mem['h0073] = 32'h200007B7;
mem['h0074] = 32'h00878793;
mem['h0075] = 32'h00F52023;
mem['h0076] = 32'h00A4A423;
mem['h0077] = 32'h00400513;
mem['h0078] = 32'hEF9FF0EF;
mem['h0079] = 32'h200007B7;
mem['h007A] = 32'h00C78793;
mem['h007B] = 32'h00F52023;
mem['h007C] = 32'h00A4A623;
mem['h007D] = 32'h00942023;
mem['h007E] = 32'h00400513;
mem['h007F] = 32'hEDDFF0EF;
mem['h0080] = 32'h200007B7;
mem['h0081] = 32'h01078793;
mem['h0082] = 32'h00F52023;
mem['h0083] = 32'h00A42223;
mem['h0084] = 32'h00400513;
mem['h0085] = 32'hEC5FF0EF;
mem['h0086] = 32'h200007B7;
mem['h0087] = 32'h01478793;
mem['h0088] = 32'h00F52023;
mem['h0089] = 32'h00A42423;
mem['h008A] = 32'h00400513;
mem['h008B] = 32'hEADFF0EF;
mem['h008C] = 32'h200007B7;
mem['h008D] = 32'h01878793;
mem['h008E] = 32'h00F52023;
mem['h008F] = 32'h00A42623;
mem['h0090] = 32'h00400513;
mem['h0091] = 32'hE95FF0EF;
mem['h0092] = 32'h200007B7;
mem['h0093] = 32'h01C78793;
mem['h0094] = 32'h00F52023;
mem['h0095] = 32'h00A42823;
mem['h0096] = 32'h00400513;
mem['h0097] = 32'hE7DFF0EF;
mem['h0098] = 32'h200007B7;
mem['h0099] = 32'h02078793;
mem['h009A] = 32'h00F52023;
mem['h009B] = 32'h00442783;
mem['h009C] = 32'h00A42A23;
mem['h009D] = 32'h0007A703;
mem['h009E] = 32'h56800593;
mem['h009F] = 32'h00040513;
mem['h00A0] = 32'h00072783;
mem['h00A1] = 32'h100019B7;
mem['h00A2] = 32'h2007E793;
mem['h00A3] = 32'h00F72023;
mem['h00A4] = 32'hE0DFF0EF;
mem['h00A5] = 32'h59800593;
mem['h00A6] = 32'h00040513;
mem['h00A7] = 32'hE01FF0EF;
mem['h00A8] = 32'h01C00913;
mem['h00A9] = 32'h70400493;
mem['h00AA] = 32'h80098993;
mem['h00AB] = 32'hFFC00A13;
mem['h00AC] = 32'h0129D7B3;
mem['h00AD] = 32'h00F7F793;
mem['h00AE] = 32'h00F487B3;
mem['h00AF] = 32'h0007C583;
mem['h00B0] = 32'h00040513;
mem['h00B1] = 32'hFFC90913;
mem['h00B2] = 32'hDADFF0EF;
mem['h00B3] = 32'hFF4912E3;
mem['h00B4] = 32'h5AC00593;
mem['h00B5] = 32'h00040513;
mem['h00B6] = 32'hDC5FF0EF;
mem['h00B7] = 32'h00400A13;
mem['h00B8] = 32'h3E800913;
mem['h00B9] = 32'h000019B7;
mem['h00BA] = 32'h00090593;
mem['h00BB] = 32'h00098513;
mem['h00BC] = 32'h1CC000EF;
mem['h00BD] = 32'h03050593;
mem['h00BE] = 32'h0FF5F593;
mem['h00BF] = 32'h00040513;
mem['h00C0] = 32'hD75FF0EF;
mem['h00C1] = 32'h00090593;
mem['h00C2] = 32'h00098513;
mem['h00C3] = 32'h1F8000EF;
mem['h00C4] = 32'h01051993;
mem['h00C5] = 32'h00A00593;
mem['h00C6] = 32'h00090513;
mem['h00C7] = 32'h1A0000EF;
mem['h00C8] = 32'h01051913;
mem['h00C9] = 32'hFFFA0A13;
mem['h00CA] = 32'h0109D993;
mem['h00CB] = 32'h01095913;
mem['h00CC] = 32'hFA0A1CE3;
mem['h00CD] = 32'h5BC00593;
mem['h00CE] = 32'h00040513;
mem['h00CF] = 32'hD61FF0EF;
mem['h00D0] = 32'h5C800593;
mem['h00D1] = 32'h00040513;
mem['h00D2] = 32'hD55FF0EF;
mem['h00D3] = 32'h5F400D13;
mem['h00D4] = 32'h60800D93;
mem['h00D5] = 32'h61C00793;
mem['h00D6] = 32'h00F12223;
mem['h00D7] = 32'h63C00793;
mem['h00D8] = 32'h00F12423;
mem['h00D9] = 32'h800009B7;
mem['h00DA] = 32'h65400793;
mem['h00DB] = 32'hFFF98A13;
mem['h00DC] = 32'h00F12623;
mem['h00DD] = 32'h00100713;
mem['h00DE] = 32'h00442783;
mem['h00DF] = 32'h0007A783;
mem['h00E0] = 32'h0007A783;
mem['h00E1] = 32'h0017F793;
mem['h00E2] = 32'hFEE798E3;
mem['h00E3] = 32'h000D0593;
mem['h00E4] = 32'h00040513;
mem['h00E5] = 32'hD09FF0EF;
mem['h00E6] = 32'h000D8593;
mem['h00E7] = 32'h00040513;
mem['h00E8] = 32'hCFDFF0EF;
mem['h00E9] = 32'h00C42783;
mem['h00EA] = 32'h00412583;
mem['h00EB] = 32'h00040513;
mem['h00EC] = 32'h0007A703;
mem['h00ED] = 32'h00072783;
mem['h00EE] = 32'h0137E7B3;
mem['h00EF] = 32'h00F72023;
mem['h00F0] = 32'h00C42783;
mem['h00F1] = 32'h0007A703;
mem['h00F2] = 32'h00072783;
mem['h00F3] = 32'h0147F7B3;
mem['h00F4] = 32'h00F72023;
mem['h00F5] = 32'hCC9FF0EF;
mem['h00F6] = 32'h00812583;
mem['h00F7] = 32'h00040513;
mem['h00F8] = 32'hCBDFF0EF;
mem['h00F9] = 32'h00C42783;
mem['h00FA] = 32'h0007A783;
mem['h00FB] = 32'h0007A783;
mem['h00FC] = 32'h00179713;
mem['h00FD] = 32'h0A075863;
mem['h00FE] = 32'h00C12583;
mem['h00FF] = 32'h00040513;
mem['h0100] = 32'h10001B37;
mem['h0101] = 32'hC99FF0EF;
mem['h0102] = 32'h68000593;
mem['h0103] = 32'h00040513;
mem['h0104] = 32'hC8DFF0EF;
mem['h0105] = 32'h10005937;
mem['h0106] = 32'h800B0B13;
mem['h0107] = 32'hFFC00A93;
mem['h0108] = 32'h59400C93;
mem['h0109] = 32'h80090913;
mem['h010A] = 32'h000B2C03;
mem['h010B] = 32'h01C00B93;
mem['h010C] = 32'h017C57B3;
mem['h010D] = 32'h00F7F793;
mem['h010E] = 32'h00F487B3;
mem['h010F] = 32'h0007C583;
mem['h0110] = 32'h00040513;
mem['h0111] = 32'hFFCB8B93;
mem['h0112] = 32'hC2DFF0EF;
mem['h0113] = 32'hFF5B92E3;
mem['h0114] = 32'h000C8593;
mem['h0115] = 32'h00040513;
mem['h0116] = 32'h004B0B13;
mem['h0117] = 32'hC41FF0EF;
mem['h0118] = 32'hFD2B14E3;
mem['h0119] = 32'h6A000593;
mem['h011A] = 32'h00040513;
mem['h011B] = 32'hC31FF0EF;
mem['h011C] = 32'h6BC00593;
mem['h011D] = 32'h00040513;
mem['h011E] = 32'hC25FF0EF;
mem['h011F] = 32'h6D800593;
mem['h0120] = 32'h00040513;
mem['h0121] = 32'hC19FF0EF;
mem['h0122] = 32'h00100713;
mem['h0123] = 32'h00442783;
mem['h0124] = 32'h0007A783;
mem['h0125] = 32'h0007A783;
mem['h0126] = 32'h0017F793;
mem['h0127] = 32'hECE79CE3;
mem['h0128] = 32'hFEDFF06F;
mem['h0129] = 32'h02E00593;
mem['h012A] = 32'h00040513;
mem['h012B] = 32'hBC9FF0EF;
mem['h012C] = 32'hF35FF06F;
mem['h012D] = 32'h06054063;
mem['h012E] = 32'h0605C663;
mem['h012F] = 32'h00058613;
mem['h0130] = 32'h00050593;
mem['h0131] = 32'hFFF00513;
mem['h0132] = 32'h02060C63;
mem['h0133] = 32'h00100693;
mem['h0134] = 32'h00B67A63;
mem['h0135] = 32'h00C05863;
mem['h0136] = 32'h00161613;
mem['h0137] = 32'h00169693;
mem['h0138] = 32'hFEB66AE3;
mem['h0139] = 32'h00000513;
mem['h013A] = 32'h00C5E663;
mem['h013B] = 32'h40C585B3;
mem['h013C] = 32'h00D56533;
mem['h013D] = 32'h0016D693;
mem['h013E] = 32'h00165613;
mem['h013F] = 32'hFE0696E3;
mem['h0140] = 32'h00008067;
mem['h0141] = 32'h00008293;
mem['h0142] = 32'hFB5FF0EF;
mem['h0143] = 32'h00058513;
mem['h0144] = 32'h00028067;
mem['h0145] = 32'h40A00533;
mem['h0146] = 32'h00B04863;
mem['h0147] = 32'h40B005B3;
mem['h0148] = 32'hF9DFF06F;
mem['h0149] = 32'h40B005B3;
mem['h014A] = 32'h00008293;
mem['h014B] = 32'hF91FF0EF;
mem['h014C] = 32'h40A00533;
mem['h014D] = 32'h00028067;
mem['h014E] = 32'h00008293;
mem['h014F] = 32'h0005CA63;
mem['h0150] = 32'h00054C63;
mem['h0151] = 32'hF79FF0EF;
mem['h0152] = 32'h00058513;
mem['h0153] = 32'h00028067;
mem['h0154] = 32'h40B005B3;
mem['h0155] = 32'hFE0558E3;
mem['h0156] = 32'h40A00533;
mem['h0157] = 32'hF61FF0EF;
mem['h0158] = 32'h40B00533;
mem['h0159] = 32'h00028067;
mem['h015A] = 32'h202D2D2D;
mem['h015B] = 32'h43534952;
mem['h015C] = 32'h4120562D;
mem['h015D] = 32'h53204344;
mem['h015E] = 32'h7370616E;
mem['h015F] = 32'h20746F68;
mem['h0160] = 32'h75716341;
mem['h0161] = 32'h74697369;
mem['h0162] = 32'h206E6F69;
mem['h0163] = 32'h6F6D6544;
mem['h0164] = 32'h2D2D2D20;
mem['h0165] = 32'h00000A0D;
mem['h0166] = 32'h66667542;
mem['h0167] = 32'h61207265;
mem['h0168] = 32'h73657264;
mem['h0169] = 32'h30203A61;
mem['h016A] = 32'h00000078;
mem['h016B] = 32'h6556202C;
mem['h016C] = 32'h6963696C;
mem['h016D] = 32'h203A616E;
mem['h016E] = 32'h00000000;
mem['h016F] = 32'h6F7A7520;
mem['h0170] = 32'h616B6172;
mem['h0171] = 32'h000A0D2E;
mem['h0172] = 32'h74697250;
mem['h0173] = 32'h696E7369;
mem['h0174] = 32'h4B206574;
mem['h0175] = 32'h20315945;
mem['h0176] = 32'h4620616E;
mem['h0177] = 32'h20414750;
mem['h0178] = 32'h6120617A;
mem['h0179] = 32'h7A69766B;
mem['h017A] = 32'h6A696369;
mem['h017B] = 32'h2E2E2E75;
mem['h017C] = 32'h00000A0D;
mem['h017D] = 32'h74697250;
mem['h017E] = 32'h756E7369;
mem['h017F] = 32'h454B2074;
mem['h0180] = 32'h0D2E3159;
mem['h0181] = 32'h0000000A;
mem['h0182] = 32'h3A434441;
mem['h0183] = 32'h69725020;
mem['h0184] = 32'h6D657270;
mem['h0185] = 32'h2E2E2E61;
mem['h0186] = 32'h00000A0D;
mem['h0187] = 32'h3A434441;
mem['h0188] = 32'h766B4120;
mem['h0189] = 32'h63697A69;
mem['h018A] = 32'h20616A69;
mem['h018B] = 32'h6F70617A;
mem['h018C] = 32'h61746563;
mem['h018D] = 32'h0D2E2E2E;
mem['h018E] = 32'h0000000A;
mem['h018F] = 32'h3A434441;
mem['h0190] = 32'h6B654320;
mem['h0191] = 32'h206F6D61;
mem['h0192] = 32'h656E6F64;
mem['h0193] = 32'h0D2E2E2E;
mem['h0194] = 32'h0000000A;
mem['h0195] = 32'h3A434441;
mem['h0196] = 32'h66614220;
mem['h0197] = 32'h70207265;
mem['h0198] = 32'h6E75706F;
mem['h0199] = 32'h2E6E656A;
mem['h019A] = 32'h6B6F5020;
mem['h019B] = 32'h65636572;
mem['h019C] = 32'h7274206D;
mem['h019D] = 32'h66736E61;
mem['h019E] = 32'h2E2E7265;
mem['h019F] = 32'h000A0D2E;
mem['h01A0] = 32'h203D3D3D;
mem['h01A1] = 32'h4D415242;
mem['h01A2] = 32'h4152545F;
mem['h01A3] = 32'h4546534E;
mem['h01A4] = 32'h54535F52;
mem['h01A5] = 32'h20545241;
mem['h01A6] = 32'h0D3D3D3D;
mem['h01A7] = 32'h0000000A;
mem['h01A8] = 32'h203D3D3D;
mem['h01A9] = 32'h4D415242;
mem['h01AA] = 32'h4152545F;
mem['h01AB] = 32'h4546534E;
mem['h01AC] = 32'h4E455F52;
mem['h01AD] = 32'h3D3D2044;
mem['h01AE] = 32'h000A0D3D;
mem['h01AF] = 32'h3A434441;
mem['h01B0] = 32'h61725420;
mem['h01B1] = 32'h6566736E;
mem['h01B2] = 32'h617A2072;
mem['h01B3] = 32'h65737276;
mem['h01B4] = 32'h0A0D2E6E;
mem['h01B5] = 32'h00000000;
mem['h01B6] = 32'h65727053;
mem['h01B7] = 32'h206E616D;
mem['h01B8] = 32'h6E20617A;
mem['h01B9] = 32'h2075766F;
mem['h01BA] = 32'h69766B61;
mem['h01BB] = 32'h6963697A;
mem['h01BC] = 32'h2820756A;
mem['h01BD] = 32'h616B6543;
mem['h01BE] = 32'h454B206D;
mem['h01BF] = 32'h2E293159;
mem['h01C0] = 32'h00000A0D;
mem['h01C1] = 32'h33323130;
mem['h01C2] = 32'h37363534;
mem['h01C3] = 32'h42413938;
mem['h01C4] = 32'h46454443;
mem['h01C5] = 32'h00000000;
